// Tasks file for producing instructions.

task rtype_insn (
  input logic [6:0] opcode,
  input logic [4:0] rd,
  input logic [2:0] funct3,
  input [4:0] rs1,
  input [4:0] rs2,
  input [6:0] funct7,
  output [31:0] insn
);
  begin
    insn = {funct7, rs2, rs1, funct3, rd, opcode};
  end
endtask


task itype_insn (
  input [6:0] opcode,
  input [4:0] rd,
  input [2:0] funct3,
  input [4:0] rs1,
  input [11:0] imm,
  output [31:0] insn
);
  begin
    insn = {imm, rs1, funct3, rd, opcode};
  end
endtask

task stype_insn (
  input [6:0] opcode,
  input [2:0] funct3,
  input [4:0] rs1,
  input [4:0] rs2,
  input [11:0] imm,
  output [31:0] insn
);
  begin
    insn = {imm[11:5], rs2[4:0], rs1[4:0], funct3[2:0], imm[4:0], opcode[6:0]};
  end
endtask

task btype_insn (
  input [6:0] opcode,
  input [2:0] funct3,
  input [4:0] rs1,
  input [4:0] rs2,
  input [12:0] imm,
  output [31:0] insn
);
  begin
    insn = {imm[12], imm[10:5], rs2[4:0], rs1[4:0], funct3[2:0], imm[4:1], imm[11], opcode[6:0]};
  end
endtask

task utype_insn (
  input [6:0] opcode,
  input [4:0] rd,
  input [19:0] imm,
  output [31:0] insn
);
  begin
    insn = {imm, rd, opcode};
  end
endtask

task jtype_insn (
  input [6:0] opcode,
  input [4:0] rd,
  input [19:0] imm,
  output [31:0] insn
);
  begin
    insn = {imm[20], imm[10:1], imm[11], imm[19:12], rd[4:0], opcode[6:0]};
  end
endtask
