// ----  Probes  ----
`define PROBE_ADDR memory_addr_i      
`define PROBE_DATA_IN memory_data_i
`define PROBE_DATA_OUT insn_o  
`define PROBE_READ_EN memory_read_en_i
`define PROBE_WRITE_EN memory_write_en_i
`define PROBE_VALID   memory_valid_o

`define PROBE_F_PC fetch_pc_o
`define PROBE_F_INSN insn_o
// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd1
// ----  Top module  ----
